module test_sample();

// Declare inputs as regs and outputs as wires
reg clock;
reg init;

wire [7:0] alu_result;
wire [7:0] pc_out;
//wire mem_write_ctrl;
//wire mem_read_ctrl;
//wire [8:0] instruction;
wire [16:0] cycle_count;

// Initialize all variables
initial begin

	clock = 1; 		// initial value of clock
	
	/* 
	 * Check the sum operation 
	 */
	#10 
	//register_one = 8'b11;	// r1 = 3
	//register_two = 8'b10;		// r2 = 2
	//function_control = 4'b0;	// sum (3 + 2) = 5
	
	#10;
	//register_one = 8'b1111_1101;	// r1 = -3
	//register_two = 8'b1111_1101;	// r2 = -3
	#10;
	#10;
	#10;
	#10;
	#10;
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
	
end

// Clock generator
always begin
	#5 clock = ~clock; // Toggle clock every 5 ticks
	// this makes the clock cycle 10 ticks
end

// I copied this code verbatim from the alu_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
wire	[8:0] instruction;
wire	mem_read;
wire	SYNTHESIZED_WIRE_0;
wire	[7:0] SYNTHESIZED_WIRE_25;
wire	[7:0] SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	[3:0] SYNTHESIZED_WIRE_5;
wire	[7:0] SYNTHESIZED_WIRE_7;
wire	[2:0] SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	[1:0] SYNTHESIZED_WIRE_12;
wire	[2:0] SYNTHESIZED_WIRE_13;
wire	[7:0] SYNTHESIZED_WIRE_14;
wire	[7:0] SYNTHESIZED_WIRE_15;
wire	[7:0] SYNTHESIZED_WIRE_16;
wire	[7:0] SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	[7:0] SYNTHESIZED_WIRE_23;

assign	alu_result = SYNTHESIZED_WIRE_15;
assign	pc_out = SYNTHESIZED_WIRE_17;




control_unit	b2v_inst(
	.clock(clock),
	.instruction(instruction),
	.alu_src(SYNTHESIZED_WIRE_18),
	.mem_write(SYNTHESIZED_WIRE_0),
	.mem_read(mem_read),
	.branch(SYNTHESIZED_WIRE_3),
	.reg_write(SYNTHESIZED_WIRE_9),
	.swap_ctrl(SYNTHESIZED_WIRE_11),
	.done_ctrl(SYNTHESIZED_WIRE_22),
	.jmp_ctrl(SYNTHESIZED_WIRE_21),
	.alu_func(SYNTHESIZED_WIRE_5),
	.alu_spec_func(SYNTHESIZED_WIRE_8),
	.reg_write_val(SYNTHESIZED_WIRE_13),
	.set_ctrl(SYNTHESIZED_WIRE_12));


single_port_ram_with_init	b2v_inst1(
	.writemem(SYNTHESIZED_WIRE_0),
	.readmem(mem_read),
	.clk(clock),
	.addr(SYNTHESIZED_WIRE_25),
	.data(SYNTHESIZED_WIRE_26),
	.q(SYNTHESIZED_WIRE_16));
	defparam	b2v_inst1.ADDR_WIDTH = 8;

assign	SYNTHESIZED_WIRE_20 = SYNTHESIZED_WIRE_3 & SYNTHESIZED_WIRE_4;


alu	b2v_inst4(
	.clock(clock),
	.func(SYNTHESIZED_WIRE_5),
	.reg1(SYNTHESIZED_WIRE_26),
	.reg2(SYNTHESIZED_WIRE_7),
	.spec_fun(SYNTHESIZED_WIRE_8),
	.carry_out(SYNTHESIZED_WIRE_10),
	.br_out(SYNTHESIZED_WIRE_4),
	.res(SYNTHESIZED_WIRE_15));


register_file	b2v_inst5(
	.clock(clock),
	.write_ctrl(SYNTHESIZED_WIRE_9),
	.carry_out(SYNTHESIZED_WIRE_10),
	.swap_ctrl(SYNTHESIZED_WIRE_11),
	.read_reg1(instruction[4:3]),
	.read_reg2(instruction[2:0]),
	.set_ctrl(SYNTHESIZED_WIRE_12),
	.write_reg(SYNTHESIZED_WIRE_13),
	.write_val(SYNTHESIZED_WIRE_14),
	.branch_val(SYNTHESIZED_WIRE_23),
	.read_val1(SYNTHESIZED_WIRE_26),
	.read_val2(SYNTHESIZED_WIRE_25));


mux_reg_write_val	b2v_inst6(
	.selector(mem_read),
	.alu_result(SYNTHESIZED_WIRE_15),
	.mem_val(SYNTHESIZED_WIRE_16),
	.mux_reg_out(SYNTHESIZED_WIRE_14));


Instruction_rom_sample	b2v_inst7(
	.address(SYNTHESIZED_WIRE_17),
	.instruction(instruction));


mux_alu	b2v_inst8(
	.selector(SYNTHESIZED_WIRE_18),
	.immediate(instruction[3:0]),
	.register_2(SYNTHESIZED_WIRE_25),
	.mux_alu_out(SYNTHESIZED_WIRE_7));


fetch_unit	b2v_inst9(
	.clock(clock),
	.branch_ctrl(SYNTHESIZED_WIRE_20),
	.jump_ctrl(SYNTHESIZED_WIRE_21),
	.done_ctrl(SYNTHESIZED_WIRE_22),
	.init_ctrl(init),
	.branch_val(SYNTHESIZED_WIRE_23),
	.jump_val(SYNTHESIZED_WIRE_26),
	.cycle_counter(cycle_count),
	.instruction_number(SYNTHESIZED_WIRE_17));


endmodule
