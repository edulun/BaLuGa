module test_sample();

// Declare inputs as regs and outputs as wires
reg clock;
reg init;

wire [7:0] alu_result;
wire [7:0] pc_out;
wire mem_write_ctrl;
wire mem_read_ctrl;
//wire [8:0] instruction;
wire [16:0] cycle_count;

// Initialize all variables
initial begin

	clock = 1; 		// initial value of clock
	
	/* 
	 * Check the sum operation 
	 */
	#10 
	//register_one = 8'b11;	// r1 = 3
	//register_two = 8'b10;		// r2 = 2
	//function_control = 4'b0;	// sum (3 + 2) = 5
	
	#10;
	//register_one = 8'b1111_1101;	// r1 = -3
	//register_two = 8'b1111_1101;	// r2 = -3
	#10;
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
    #10;// sum (-3 + -3) = -6
	
end

// Clock generator
always begin
	#5 clock = ~clock; // Toggle clock every 5 ticks
	// this makes the clock cycle 10 ticks
end

// I copied this code verbatim from the alu_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
wire	[8:0] instruction;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	[3:0] SYNTHESIZED_WIRE_2;
wire	[7:0] SYNTHESIZED_WIRE_20;
wire	[7:0] SYNTHESIZED_WIRE_4;
wire	[2:0] SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	[1:0] SYNTHESIZED_WIRE_9;
wire	[2:0] SYNTHESIZED_WIRE_10;
wire	[7:0] SYNTHESIZED_WIRE_11;
wire	[7:0] SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	[7:0] SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	[7:0] SYNTHESIZED_WIRE_18;

assign	alu_result = SYNTHESIZED_WIRE_11;
assign	pc_out = SYNTHESIZED_WIRE_12;




control_unit	b2v_inst(
	.clock(clock),
	.instruction(instruction),
	.alu_src(SYNTHESIZED_WIRE_13),
	.mem_write(mem_write_ctrl),
	.mem_read(mem_read_ctrl),
	.branch(SYNTHESIZED_WIRE_0),
	.reg_write(SYNTHESIZED_WIRE_6),
	.swap_ctrl(SYNTHESIZED_WIRE_8),
	.done_ctrl(SYNTHESIZED_WIRE_17),
	.jmp_ctrl(SYNTHESIZED_WIRE_16),
	.alu_func(SYNTHESIZED_WIRE_2),
	.alu_spec_func(SYNTHESIZED_WIRE_5),
	.reg_write_val(SYNTHESIZED_WIRE_10),
	.set_ctrl(SYNTHESIZED_WIRE_9));

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_0 & SYNTHESIZED_WIRE_1;


alu	b2v_inst4(
	.clock(clock),
	.func(SYNTHESIZED_WIRE_2),
	.reg1(SYNTHESIZED_WIRE_20),
	.reg2(SYNTHESIZED_WIRE_4),
	.spec_fun(SYNTHESIZED_WIRE_5),
	.carry_out(SYNTHESIZED_WIRE_7),
	.br_out(SYNTHESIZED_WIRE_1),
	.res(SYNTHESIZED_WIRE_11));


register_file	b2v_inst5(
	.clock(clock),
	.write_ctrl(SYNTHESIZED_WIRE_6),
	.carry_out(SYNTHESIZED_WIRE_7),
	.swap_ctrl(SYNTHESIZED_WIRE_8),
	.read_reg1(instruction[4:3]),
	.read_reg2(instruction[2:0]),
	.set_ctrl(SYNTHESIZED_WIRE_9),
	.write_reg(SYNTHESIZED_WIRE_10),
	.write_val(SYNTHESIZED_WIRE_11),
	.branch_val(SYNTHESIZED_WIRE_18),
	.read_val1(SYNTHESIZED_WIRE_20),
	.read_val2(SYNTHESIZED_WIRE_14));


Instruction_rom_sample	b2v_inst7(
	.address(SYNTHESIZED_WIRE_12),
	.instruction(instruction));


mux_alu	b2v_inst8(
	.selector(SYNTHESIZED_WIRE_13),
	.immediate(instruction[3:0]),
	.register_2(SYNTHESIZED_WIRE_14),
	.mux_alu_out(SYNTHESIZED_WIRE_4));


fetch_unit	b2v_inst9(
	.clock(clock),
	.branch_ctrl(SYNTHESIZED_WIRE_15),
	.jump_ctrl(SYNTHESIZED_WIRE_16),
	.done_ctrl(SYNTHESIZED_WIRE_17),
	.init_ctrl(init),
	.branch_val(SYNTHESIZED_WIRE_18),
	.jump_val(SYNTHESIZED_WIRE_20),
	.cycle_counter(cycle_count),
	.instruction_number(SYNTHESIZED_WIRE_12));

endmodule
