module testbench_regFile();

// Declare inputs as regs and outputs as wires
reg clock;
reg write_ctrl;
reg swap_ctrl;
reg [1:0] read_reg1;
reg [2:0] read_reg2;
reg [2:0] write_reg;
reg [7:0] write_val;

wire [7:0] read_val1;
wire [7:0] read_val2;

// Initialize all variables
initial begin

	clock = 1; 		// initial value of clock
	write_ctrl = 0;
	swap_ctrl = 0;
	
	// 10 PS
	// Write values to regs
	// No output to read_regs
	#10 write_val = 8'd1; write_reg = 3'd1;  write_ctrl = 1; // imm = 1
	#10 write_val = 8'd2; write_reg = 3'd2;  write_ctrl = 1; // t1 = 2
	#10 write_val = 8'd3; write_reg = 3'd3;  write_ctrl = 1; // t2 = 3
	#10 write_val = 8'd4; write_reg = 3'd4;  write_ctrl = 1; // s1 = 4
	#10 write_val = 8'd5; write_reg = 3'd5;  write_ctrl = 1; // s2 = 5
	#10 write_val = 8'd6; write_reg = 3'd6;  write_ctrl = 1; // s3 = 6
	#10 write_val = 8'd7; write_reg = 3'd7;  write_ctrl = 1; // branch = 7
	
	// 80 PS
	// Read values from regs
	#10 read_reg1 = 2'd0;	read_reg2 = 3'd4;  write_ctrl = 0; //read_val1 = 0[zero], read_val1 = 4[s1]
	#10 read_reg1 = 2'd1;	read_reg2 = 3'd5;  write_ctrl = 0; //read_val1 = 1[imm], :w
	#10 read_reg1 = 2'd2;	read_reg2 = 3'd6;  write_ctrl = 0; //t1 && s3
	#10 read_reg1 = 2'd3;	read_reg2 = 3'd7;  write_ctrl = 0; //t2 && br
	#10 swap_ctrl = 1; 	read_reg1 = 2'd1;  read_reg2 = 3'd4;	  //swap imm <> s1
	
	#10 swap_ctrl = 0;
	
end

// Clock generator
always begin
	#5 clock = ~clock; // Toggle clock every 5 ticks
	// this makes the clock cycle 10 ticks
end

// I copied this code verbatim from the alu_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
register_file	b2v_inst(
	.clock(clock),
	.write_ctrl(write_ctrl),
	.swap_ctrl(swap_ctrl),
	.read_reg1(read_reg1),
	.read_reg2(read_reg2),
	.write_reg(write_reg),
	.write_val(write_val),
	.reg_val1(reg_val1),
	.reg_val2(reg_val2));




endmodule
