module testbench_regFile();

// Declare inputs as regs and outputs as wires
reg clock;
reg wrCtrl;
reg swapCtrl;
reg [1:0] reg1;
reg [2:0] reg2;
reg [2:0] wr_reg;
reg [7:0] wr_data;

wire [7:0] regVal1;
wire [7:0] regVal2;

// Initialize all variables
initial begin

	clock = 1; 		// initial value of clock
	wrCtrl = 0;
	swapCtrl = 0;
	
	
	#10 wr_data = 8'b01010101; wr_reg = 3'b010;  wrCtrl = 1;
	#10 wrCtrl = 0; wr_data = 8'b00000000;	//Register 010 shouldn't change
	#10 wr_data = 8'b00000001; wr_reg = 3'b001;  wrCtrl = 1;
	#10 wr_data = 8'b00000010; wr_reg = 3'b010;  wrCtrl = 1;
	#10 wr_data = 8'b00000011; wr_reg = 3'b011;  wrCtrl = 1;
	#10 wr_data = 8'b00000100; wr_reg = 3'b100;  wrCtrl = 1;
	#10 wr_data = 8'b00000101; wr_reg = 3'b101;  wrCtrl = 1;
	#10 wr_data = 8'b00000110; wr_reg = 3'b110;  wrCtrl = 1;
	#10 wrCtrl = 0;
	#10 reg1 = 2'b00; reg2 = 3'b001;
	#10 reg1 = 2'b11; reg2 = 3'b101; swapCtrl = 1;
	#10 swapCtrl = 0;
end

// Clock generator
always begin
	#5 clock = ~clock; // Toggle clock every 5 ticks
	// this makes the clock cycle 10 ticks
end

// I copied this code verbatim from the alu_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
register_file	b2v_inst(
	.clock(clock),
	.write_to_reg(wrCtrl),
	.swap_regs(swapCtrl),
	.rd_reg1(reg1),
	.rd_reg2(reg2),
	.wr_reg(wr_reg),
	.write_data(wr_data),
	.reg_val1(regVal1),
	.reg_val2(regVal2));

endmodule