module test_bench_control_unit();

// Declare inputs as regs and outputs as wires
reg clock;
reg [8:0] instr;

wire [6:0] alu_ctrl;
wire [2:0] reg_to_write;
wire alu_mux_ctrl;
wire mem_write;
wire mem_read;
wire branch;
wire reg_write;
wire swap_ctrl;
wire done_ctrl;
wire jump_ctrl;

// Initialize all variables
initial begin

	clock = 1; 		// initial value of clock
	
	/* 
	 * Check the sum instruction 
	 */
	#10; 
	instr = 9'b0000_10_100;		// add $2,$4
	// Expected ouput:
	// alu_ctrl = 0000XX
	// reg_to_write = 010
	// mem_write = 0
	// mem_read = 0
	// wire branch = 0
	// reg_write = 1
	// swap_ctrl = 0
	// done_ctrl = 0
	// jump_ctrl = 0 	
end

// Clock generator
always begin
	#5 clock = ~clock; // Toggle clock every 5 ticks
	// this makes the clock cycle 10 ticks
end

// I copied this code verbatim from the alu_schematic.v that was
// generated by Quartus when I created the .v file from the .bdf.
control_unit	b2v_inst(
	.clock(clock),
	.instruction(instr),
	.alu_src(alu_mux_ctrl),
	.mem_write(mem_write),
	.mem_read(mem_read),
	.branch(branch),
	.reg_write(reg_write),
	.swap_ctrl(swap_ctrl),
	.done_ctrl(done_ctrl),
	.jmp_ctrl(jump_ctrl),
	.alu_ctrl(alu_ctrl),
	.reg_write_val(reg_to_write));


endmodule